parameter int DATA_SIZE = 8;
parameter int INST_SIZE = 16;
parameter int MEM_DEPTH = 128;
